enum { circle, ellipse, freeform } c;
